// DE0_CV_QSYS.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module DE0_CV_QSYS (
		input  wire        clk_clk,                                     //                              clk.clk
		output wire        clk_5m_clk,                                  //                           clk_5m.clk
		output wire        clk_sdram_clk,                               //                        clk_sdram.clk
		output wire        ltc2992_i2c_sda_t,                           //                      ltc2992_i2c.sda_t
		output wire        ltc2992_i2c_scl_t,                           //                                 .scl_t
		input  wire        ltc2992_i2c_sda_i,                           //                                 .sda_i
		input  wire        ltc2992_i2c_scl_i,                           //                                 .scl_i
		output wire        pll_locked_export,                           //                       pll_locked.export
		input  wire        reset_reset_n,                               //                            reset.reset_n
		output wire [12:0] sdram_wire_addr,                             //                       sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                               //                                 .ba
		output wire        sdram_wire_cas_n,                            //                                 .cas_n
		output wire        sdram_wire_cke,                              //                                 .cke
		output wire        sdram_wire_cs_n,                             //                                 .cs_n
		inout  wire [15:0] sdram_wire_dq,                               //                                 .dq
		output wire [1:0]  sdram_wire_dqm,                              //                                 .dqm
		output wire        sdram_wire_ras_n,                            //                                 .ras_n
		output wire        sdram_wire_we_n,                             //                                 .we_n
		output wire        servo_controllerv1_0_conduit_end_spi_sclk,   // servo_controllerv1_0_conduit_end.spi_sclk
		output wire        servo_controllerv1_0_conduit_end_spi_cs,     //                                 .spi_cs
		input  wire        servo_controllerv1_0_conduit_end_spi_miso,   //                                 .spi_miso
		output wire        servo_controllerv1_0_conduit_end_spi_mosi,   //                                 .spi_mosi
		input  wire [2:0]  servo_controllerv1_0_conduit_end_hall_0,     //                                 .hall_0
		input  wire [2:0]  servo_controllerv1_0_conduit_end_hall_1,     //                                 .hall_1
		input  wire [2:0]  servo_controllerv1_0_conduit_end_hall_2,     //                                 .hall_2
		input  wire [2:0]  servo_controllerv1_0_conduit_end_hall_3,     //                                 .hall_3
		output wire [5:0]  servo_controllerv1_0_conduit_end_phase_0,    //                                 .phase_0
		output wire [5:0]  servo_controllerv1_0_conduit_end_phase_1,    //                                 .phase_1
		output wire [5:0]  servo_controllerv1_0_conduit_end_phase_2,    //                                 .phase_2
		output wire [5:0]  servo_controllerv1_0_conduit_end_phase_3,    //                                 .phase_3
		input  wire [3:0]  servo_controllerv1_0_conduit_end_nFault,     //                                 .nFault
		output wire [3:0]  servo_controllerv1_0_conduit_end_drv8320_en, //                                 .drv8320_en
		output wire        tmp101_i2c_sda_t,                            //                       tmp101_i2c.sda_t
		output wire        tmp101_i2c_scl_t,                            //                                 .scl_t
		input  wire        tmp101_i2c_sda_i,                            //                                 .sda_i
		input  wire        tmp101_i2c_scl_i,                            //                                 .scl_i
		input  wire        uart_rs485_conduit_end_rxd,                  //           uart_rs485_conduit_end.rxd
		output wire        uart_rs485_conduit_end_txd,                  //                                 .txd
		output wire        uart_rs485_conduit_end_dbg_os_pulse          //                                 .dbg_os_pulse
	);

	wire         pll_outclk0_clk;                                                                  // pll:outclk_0 -> [boot_rom:clk, boot_rom:clk2, epcs_flash_controller_0:clk, irq_mapper:clk, jtag_uart:clk, ltc2992:clk, mm_interconnect_0:pll_outclk0_clk, mm_interconnect_1:pll_outclk0_clk, mm_interconnect_2:pll_outclk0_clk, nios2_qsys:clk, rst_controller:clk, rst_controller_001:clk, sdram:clk, servo_controllerv1_0:clk, sysid_qsys:clock, tc_instruct_mem:clk, tc_instruct_mem:clk2, timer:clk, timestamp:clk, tmp101:clk, uart_rs485:clk]
	wire         nios2_qsys_custom_instruction_master_readra;                                      // nios2_qsys:E_ci_combo_readra -> nios2_qsys_custom_instruction_master_translator:ci_slave_readra
	wire         nios2_qsys_custom_instruction_master_readrb;                                      // nios2_qsys:E_ci_combo_readrb -> nios2_qsys_custom_instruction_master_translator:ci_slave_readrb
	wire   [4:0] nios2_qsys_custom_instruction_master_multi_b;                                     // nios2_qsys:A_ci_multi_b -> nios2_qsys_custom_instruction_master_translator:ci_slave_multi_b
	wire   [4:0] nios2_qsys_custom_instruction_master_multi_c;                                     // nios2_qsys:A_ci_multi_c -> nios2_qsys_custom_instruction_master_translator:ci_slave_multi_c
	wire         nios2_qsys_custom_instruction_master_reset_req;                                   // nios2_qsys:A_ci_multi_reset_req -> nios2_qsys_custom_instruction_master_translator:ci_slave_multi_reset_req
	wire   [4:0] nios2_qsys_custom_instruction_master_multi_a;                                     // nios2_qsys:A_ci_multi_a -> nios2_qsys_custom_instruction_master_translator:ci_slave_multi_a
	wire  [31:0] nios2_qsys_custom_instruction_master_result;                                      // nios2_qsys_custom_instruction_master_translator:ci_slave_result -> nios2_qsys:E_ci_combo_result
	wire  [31:0] nios2_qsys_custom_instruction_master_datab;                                       // nios2_qsys:E_ci_combo_datab -> nios2_qsys_custom_instruction_master_translator:ci_slave_datab
	wire  [31:0] nios2_qsys_custom_instruction_master_dataa;                                       // nios2_qsys:E_ci_combo_dataa -> nios2_qsys_custom_instruction_master_translator:ci_slave_dataa
	wire         nios2_qsys_custom_instruction_master_writerc;                                     // nios2_qsys:E_ci_combo_writerc -> nios2_qsys_custom_instruction_master_translator:ci_slave_writerc
	wire  [31:0] nios2_qsys_custom_instruction_master_multi_dataa;                                 // nios2_qsys:A_ci_multi_dataa -> nios2_qsys_custom_instruction_master_translator:ci_slave_multi_dataa
	wire         nios2_qsys_custom_instruction_master_multi_writerc;                               // nios2_qsys:A_ci_multi_writerc -> nios2_qsys_custom_instruction_master_translator:ci_slave_multi_writerc
	wire   [4:0] nios2_qsys_custom_instruction_master_a;                                           // nios2_qsys:E_ci_combo_a -> nios2_qsys_custom_instruction_master_translator:ci_slave_a
	wire   [4:0] nios2_qsys_custom_instruction_master_b;                                           // nios2_qsys:E_ci_combo_b -> nios2_qsys_custom_instruction_master_translator:ci_slave_b
	wire  [31:0] nios2_qsys_custom_instruction_master_multi_result;                                // nios2_qsys_custom_instruction_master_translator:ci_slave_multi_result -> nios2_qsys:A_ci_multi_result
	wire         nios2_qsys_custom_instruction_master_clk;                                         // nios2_qsys:A_ci_multi_clock -> nios2_qsys_custom_instruction_master_translator:ci_slave_multi_clk
	wire  [31:0] nios2_qsys_custom_instruction_master_multi_datab;                                 // nios2_qsys:A_ci_multi_datab -> nios2_qsys_custom_instruction_master_translator:ci_slave_multi_datab
	wire   [4:0] nios2_qsys_custom_instruction_master_c;                                           // nios2_qsys:E_ci_combo_c -> nios2_qsys_custom_instruction_master_translator:ci_slave_c
	wire  [31:0] nios2_qsys_custom_instruction_master_ipending;                                    // nios2_qsys:E_ci_combo_ipending -> nios2_qsys_custom_instruction_master_translator:ci_slave_ipending
	wire         nios2_qsys_custom_instruction_master_start;                                       // nios2_qsys:A_ci_multi_start -> nios2_qsys_custom_instruction_master_translator:ci_slave_multi_start
	wire         nios2_qsys_custom_instruction_master_done;                                        // nios2_qsys_custom_instruction_master_translator:ci_slave_multi_done -> nios2_qsys:A_ci_multi_done
	wire   [7:0] nios2_qsys_custom_instruction_master_n;                                           // nios2_qsys:E_ci_combo_n -> nios2_qsys_custom_instruction_master_translator:ci_slave_n
	wire         nios2_qsys_custom_instruction_master_estatus;                                     // nios2_qsys:E_ci_combo_estatus -> nios2_qsys_custom_instruction_master_translator:ci_slave_estatus
	wire         nios2_qsys_custom_instruction_master_clk_en;                                      // nios2_qsys:A_ci_multi_clk_en -> nios2_qsys_custom_instruction_master_translator:ci_slave_multi_clken
	wire         nios2_qsys_custom_instruction_master_reset;                                       // nios2_qsys:A_ci_multi_reset -> nios2_qsys_custom_instruction_master_translator:ci_slave_multi_reset
	wire         nios2_qsys_custom_instruction_master_multi_readrb;                                // nios2_qsys:A_ci_multi_readrb -> nios2_qsys_custom_instruction_master_translator:ci_slave_multi_readrb
	wire         nios2_qsys_custom_instruction_master_multi_readra;                                // nios2_qsys:A_ci_multi_readra -> nios2_qsys_custom_instruction_master_translator:ci_slave_multi_readra
	wire   [7:0] nios2_qsys_custom_instruction_master_multi_n;                                     // nios2_qsys:A_ci_multi_n -> nios2_qsys_custom_instruction_master_translator:ci_slave_multi_n
	wire  [31:0] nios2_qsys_custom_instruction_master_translator_comb_ci_master_result;            // nios2_qsys_custom_instruction_master_comb_xconnect:ci_slave_result -> nios2_qsys_custom_instruction_master_translator:comb_ci_master_result
	wire         nios2_qsys_custom_instruction_master_translator_comb_ci_master_readra;            // nios2_qsys_custom_instruction_master_translator:comb_ci_master_readra -> nios2_qsys_custom_instruction_master_comb_xconnect:ci_slave_readra
	wire   [4:0] nios2_qsys_custom_instruction_master_translator_comb_ci_master_a;                 // nios2_qsys_custom_instruction_master_translator:comb_ci_master_a -> nios2_qsys_custom_instruction_master_comb_xconnect:ci_slave_a
	wire   [4:0] nios2_qsys_custom_instruction_master_translator_comb_ci_master_b;                 // nios2_qsys_custom_instruction_master_translator:comb_ci_master_b -> nios2_qsys_custom_instruction_master_comb_xconnect:ci_slave_b
	wire         nios2_qsys_custom_instruction_master_translator_comb_ci_master_readrb;            // nios2_qsys_custom_instruction_master_translator:comb_ci_master_readrb -> nios2_qsys_custom_instruction_master_comb_xconnect:ci_slave_readrb
	wire   [4:0] nios2_qsys_custom_instruction_master_translator_comb_ci_master_c;                 // nios2_qsys_custom_instruction_master_translator:comb_ci_master_c -> nios2_qsys_custom_instruction_master_comb_xconnect:ci_slave_c
	wire         nios2_qsys_custom_instruction_master_translator_comb_ci_master_estatus;           // nios2_qsys_custom_instruction_master_translator:comb_ci_master_estatus -> nios2_qsys_custom_instruction_master_comb_xconnect:ci_slave_estatus
	wire  [31:0] nios2_qsys_custom_instruction_master_translator_comb_ci_master_ipending;          // nios2_qsys_custom_instruction_master_translator:comb_ci_master_ipending -> nios2_qsys_custom_instruction_master_comb_xconnect:ci_slave_ipending
	wire  [31:0] nios2_qsys_custom_instruction_master_translator_comb_ci_master_datab;             // nios2_qsys_custom_instruction_master_translator:comb_ci_master_datab -> nios2_qsys_custom_instruction_master_comb_xconnect:ci_slave_datab
	wire  [31:0] nios2_qsys_custom_instruction_master_translator_comb_ci_master_dataa;             // nios2_qsys_custom_instruction_master_translator:comb_ci_master_dataa -> nios2_qsys_custom_instruction_master_comb_xconnect:ci_slave_dataa
	wire         nios2_qsys_custom_instruction_master_translator_comb_ci_master_writerc;           // nios2_qsys_custom_instruction_master_translator:comb_ci_master_writerc -> nios2_qsys_custom_instruction_master_comb_xconnect:ci_slave_writerc
	wire   [7:0] nios2_qsys_custom_instruction_master_translator_comb_ci_master_n;                 // nios2_qsys_custom_instruction_master_translator:comb_ci_master_n -> nios2_qsys_custom_instruction_master_comb_xconnect:ci_slave_n
	wire  [31:0] nios2_qsys_custom_instruction_master_comb_xconnect_ci_master0_result;             // nios2_qsys_custom_instruction_master_comb_slave_translator0:ci_slave_result -> nios2_qsys_custom_instruction_master_comb_xconnect:ci_master0_result
	wire         nios2_qsys_custom_instruction_master_comb_xconnect_ci_master0_readra;             // nios2_qsys_custom_instruction_master_comb_xconnect:ci_master0_readra -> nios2_qsys_custom_instruction_master_comb_slave_translator0:ci_slave_readra
	wire   [4:0] nios2_qsys_custom_instruction_master_comb_xconnect_ci_master0_a;                  // nios2_qsys_custom_instruction_master_comb_xconnect:ci_master0_a -> nios2_qsys_custom_instruction_master_comb_slave_translator0:ci_slave_a
	wire   [4:0] nios2_qsys_custom_instruction_master_comb_xconnect_ci_master0_b;                  // nios2_qsys_custom_instruction_master_comb_xconnect:ci_master0_b -> nios2_qsys_custom_instruction_master_comb_slave_translator0:ci_slave_b
	wire         nios2_qsys_custom_instruction_master_comb_xconnect_ci_master0_readrb;             // nios2_qsys_custom_instruction_master_comb_xconnect:ci_master0_readrb -> nios2_qsys_custom_instruction_master_comb_slave_translator0:ci_slave_readrb
	wire   [4:0] nios2_qsys_custom_instruction_master_comb_xconnect_ci_master0_c;                  // nios2_qsys_custom_instruction_master_comb_xconnect:ci_master0_c -> nios2_qsys_custom_instruction_master_comb_slave_translator0:ci_slave_c
	wire         nios2_qsys_custom_instruction_master_comb_xconnect_ci_master0_estatus;            // nios2_qsys_custom_instruction_master_comb_xconnect:ci_master0_estatus -> nios2_qsys_custom_instruction_master_comb_slave_translator0:ci_slave_estatus
	wire  [31:0] nios2_qsys_custom_instruction_master_comb_xconnect_ci_master0_ipending;           // nios2_qsys_custom_instruction_master_comb_xconnect:ci_master0_ipending -> nios2_qsys_custom_instruction_master_comb_slave_translator0:ci_slave_ipending
	wire  [31:0] nios2_qsys_custom_instruction_master_comb_xconnect_ci_master0_datab;              // nios2_qsys_custom_instruction_master_comb_xconnect:ci_master0_datab -> nios2_qsys_custom_instruction_master_comb_slave_translator0:ci_slave_datab
	wire  [31:0] nios2_qsys_custom_instruction_master_comb_xconnect_ci_master0_dataa;              // nios2_qsys_custom_instruction_master_comb_xconnect:ci_master0_dataa -> nios2_qsys_custom_instruction_master_comb_slave_translator0:ci_slave_dataa
	wire         nios2_qsys_custom_instruction_master_comb_xconnect_ci_master0_writerc;            // nios2_qsys_custom_instruction_master_comb_xconnect:ci_master0_writerc -> nios2_qsys_custom_instruction_master_comb_slave_translator0:ci_slave_writerc
	wire   [7:0] nios2_qsys_custom_instruction_master_comb_xconnect_ci_master0_n;                  // nios2_qsys_custom_instruction_master_comb_xconnect:ci_master0_n -> nios2_qsys_custom_instruction_master_comb_slave_translator0:ci_slave_n
	wire  [31:0] nios2_qsys_custom_instruction_master_comb_slave_translator0_ci_master_result;     // nios_custom_instr_floating_point_2_0:s1_result -> nios2_qsys_custom_instruction_master_comb_slave_translator0:ci_master_result
	wire  [31:0] nios2_qsys_custom_instruction_master_comb_slave_translator0_ci_master_datab;      // nios2_qsys_custom_instruction_master_comb_slave_translator0:ci_master_datab -> nios_custom_instr_floating_point_2_0:s1_datab
	wire  [31:0] nios2_qsys_custom_instruction_master_comb_slave_translator0_ci_master_dataa;      // nios2_qsys_custom_instruction_master_comb_slave_translator0:ci_master_dataa -> nios_custom_instr_floating_point_2_0:s1_dataa
	wire   [3:0] nios2_qsys_custom_instruction_master_comb_slave_translator0_ci_master_n;          // nios2_qsys_custom_instruction_master_comb_slave_translator0:ci_master_n -> nios_custom_instr_floating_point_2_0:s1_n
	wire         nios2_qsys_custom_instruction_master_translator_multi_ci_master_readra;           // nios2_qsys_custom_instruction_master_translator:multi_ci_master_readra -> nios2_qsys_custom_instruction_master_multi_xconnect:ci_slave_readra
	wire   [4:0] nios2_qsys_custom_instruction_master_translator_multi_ci_master_a;                // nios2_qsys_custom_instruction_master_translator:multi_ci_master_a -> nios2_qsys_custom_instruction_master_multi_xconnect:ci_slave_a
	wire   [4:0] nios2_qsys_custom_instruction_master_translator_multi_ci_master_b;                // nios2_qsys_custom_instruction_master_translator:multi_ci_master_b -> nios2_qsys_custom_instruction_master_multi_xconnect:ci_slave_b
	wire         nios2_qsys_custom_instruction_master_translator_multi_ci_master_clk;              // nios2_qsys_custom_instruction_master_translator:multi_ci_master_clk -> nios2_qsys_custom_instruction_master_multi_xconnect:ci_slave_clk
	wire         nios2_qsys_custom_instruction_master_translator_multi_ci_master_readrb;           // nios2_qsys_custom_instruction_master_translator:multi_ci_master_readrb -> nios2_qsys_custom_instruction_master_multi_xconnect:ci_slave_readrb
	wire   [4:0] nios2_qsys_custom_instruction_master_translator_multi_ci_master_c;                // nios2_qsys_custom_instruction_master_translator:multi_ci_master_c -> nios2_qsys_custom_instruction_master_multi_xconnect:ci_slave_c
	wire         nios2_qsys_custom_instruction_master_translator_multi_ci_master_start;            // nios2_qsys_custom_instruction_master_translator:multi_ci_master_start -> nios2_qsys_custom_instruction_master_multi_xconnect:ci_slave_start
	wire         nios2_qsys_custom_instruction_master_translator_multi_ci_master_reset_req;        // nios2_qsys_custom_instruction_master_translator:multi_ci_master_reset_req -> nios2_qsys_custom_instruction_master_multi_xconnect:ci_slave_reset_req
	wire         nios2_qsys_custom_instruction_master_translator_multi_ci_master_done;             // nios2_qsys_custom_instruction_master_multi_xconnect:ci_slave_done -> nios2_qsys_custom_instruction_master_translator:multi_ci_master_done
	wire   [7:0] nios2_qsys_custom_instruction_master_translator_multi_ci_master_n;                // nios2_qsys_custom_instruction_master_translator:multi_ci_master_n -> nios2_qsys_custom_instruction_master_multi_xconnect:ci_slave_n
	wire  [31:0] nios2_qsys_custom_instruction_master_translator_multi_ci_master_result;           // nios2_qsys_custom_instruction_master_multi_xconnect:ci_slave_result -> nios2_qsys_custom_instruction_master_translator:multi_ci_master_result
	wire         nios2_qsys_custom_instruction_master_translator_multi_ci_master_clk_en;           // nios2_qsys_custom_instruction_master_translator:multi_ci_master_clken -> nios2_qsys_custom_instruction_master_multi_xconnect:ci_slave_clken
	wire  [31:0] nios2_qsys_custom_instruction_master_translator_multi_ci_master_datab;            // nios2_qsys_custom_instruction_master_translator:multi_ci_master_datab -> nios2_qsys_custom_instruction_master_multi_xconnect:ci_slave_datab
	wire  [31:0] nios2_qsys_custom_instruction_master_translator_multi_ci_master_dataa;            // nios2_qsys_custom_instruction_master_translator:multi_ci_master_dataa -> nios2_qsys_custom_instruction_master_multi_xconnect:ci_slave_dataa
	wire         nios2_qsys_custom_instruction_master_translator_multi_ci_master_reset;            // nios2_qsys_custom_instruction_master_translator:multi_ci_master_reset -> nios2_qsys_custom_instruction_master_multi_xconnect:ci_slave_reset
	wire         nios2_qsys_custom_instruction_master_translator_multi_ci_master_writerc;          // nios2_qsys_custom_instruction_master_translator:multi_ci_master_writerc -> nios2_qsys_custom_instruction_master_multi_xconnect:ci_slave_writerc
	wire         nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_readra;            // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master0_readra -> nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	wire   [4:0] nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_a;                 // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master0_a -> nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_slave_a
	wire   [4:0] nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_b;                 // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master0_b -> nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_slave_b
	wire         nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_readrb;            // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master0_readrb -> nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	wire   [4:0] nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_c;                 // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master0_c -> nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_slave_c
	wire         nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_clk;               // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master0_clk -> nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	wire  [31:0] nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_ipending;          // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master0_ipending -> nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	wire         nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_start;             // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master0_start -> nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_slave_start
	wire         nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_reset_req;         // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master0_reset_req -> nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_slave_reset_req
	wire         nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_done;              // nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_slave_done -> nios2_qsys_custom_instruction_master_multi_xconnect:ci_master0_done
	wire   [7:0] nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_n;                 // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master0_n -> nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_slave_n
	wire  [31:0] nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_result;            // nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_slave_result -> nios2_qsys_custom_instruction_master_multi_xconnect:ci_master0_result
	wire         nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_estatus;           // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master0_estatus -> nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	wire         nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_clk_en;            // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master0_clken -> nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	wire  [31:0] nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_datab;             // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master0_datab -> nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	wire  [31:0] nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_dataa;             // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master0_dataa -> nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	wire         nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_reset;             // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master0_reset -> nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	wire         nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_writerc;           // nios2_qsys_custom_instruction_master_multi_xconnect:ci_master0_writerc -> nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	wire  [31:0] nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_result;    // nios_custom_instr_floating_point_2_0:s2_result -> nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_master_result
	wire         nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_clk;       // nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_master_clk -> nios_custom_instr_floating_point_2_0:s2_clk
	wire         nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_clk_en;    // nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_master_clken -> nios_custom_instr_floating_point_2_0:s2_clk_en
	wire  [31:0] nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_datab;     // nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_master_datab -> nios_custom_instr_floating_point_2_0:s2_datab
	wire  [31:0] nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_dataa;     // nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> nios_custom_instr_floating_point_2_0:s2_dataa
	wire         nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_start;     // nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_master_start -> nios_custom_instr_floating_point_2_0:s2_start
	wire         nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_reset;     // nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_master_reset -> nios_custom_instr_floating_point_2_0:s2_reset
	wire         nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_reset_req; // nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_master_reset_req -> nios_custom_instr_floating_point_2_0:s2_reset_req
	wire         nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_done;      // nios_custom_instr_floating_point_2_0:s2_done -> nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_master_done
	wire   [2:0] nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_n;         // nios2_qsys_custom_instruction_master_multi_slave_translator0:ci_master_n -> nios_custom_instr_floating_point_2_0:s2_n
	wire  [31:0] nios2_qsys_data_master_readdata;                                                  // mm_interconnect_0:nios2_qsys_data_master_readdata -> nios2_qsys:d_readdata
	wire         nios2_qsys_data_master_waitrequest;                                               // mm_interconnect_0:nios2_qsys_data_master_waitrequest -> nios2_qsys:d_waitrequest
	wire         nios2_qsys_data_master_debugaccess;                                               // nios2_qsys:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_data_master_debugaccess
	wire  [27:0] nios2_qsys_data_master_address;                                                   // nios2_qsys:d_address -> mm_interconnect_0:nios2_qsys_data_master_address
	wire   [3:0] nios2_qsys_data_master_byteenable;                                                // nios2_qsys:d_byteenable -> mm_interconnect_0:nios2_qsys_data_master_byteenable
	wire         nios2_qsys_data_master_read;                                                      // nios2_qsys:d_read -> mm_interconnect_0:nios2_qsys_data_master_read
	wire         nios2_qsys_data_master_readdatavalid;                                             // mm_interconnect_0:nios2_qsys_data_master_readdatavalid -> nios2_qsys:d_readdatavalid
	wire         nios2_qsys_data_master_write;                                                     // nios2_qsys:d_write -> mm_interconnect_0:nios2_qsys_data_master_write
	wire  [31:0] nios2_qsys_data_master_writedata;                                                 // nios2_qsys:d_writedata -> mm_interconnect_0:nios2_qsys_data_master_writedata
	wire  [31:0] nios2_qsys_instruction_master_readdata;                                           // mm_interconnect_0:nios2_qsys_instruction_master_readdata -> nios2_qsys:i_readdata
	wire         nios2_qsys_instruction_master_waitrequest;                                        // mm_interconnect_0:nios2_qsys_instruction_master_waitrequest -> nios2_qsys:i_waitrequest
	wire  [27:0] nios2_qsys_instruction_master_address;                                            // nios2_qsys:i_address -> mm_interconnect_0:nios2_qsys_instruction_master_address
	wire         nios2_qsys_instruction_master_read;                                               // nios2_qsys:i_read -> mm_interconnect_0:nios2_qsys_instruction_master_read
	wire         nios2_qsys_instruction_master_readdatavalid;                                      // mm_interconnect_0:nios2_qsys_instruction_master_readdatavalid -> nios2_qsys:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;                         // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;                           // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;                        // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;                            // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                               // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;                              // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;                          // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_servo_controllerv1_0_avalon_slave_0_readdata;                   // servo_controllerv1_0:readdata -> mm_interconnect_0:servo_controllerv1_0_avalon_slave_0_readdata
	wire   [4:0] mm_interconnect_0_servo_controllerv1_0_avalon_slave_0_address;                    // mm_interconnect_0:servo_controllerv1_0_avalon_slave_0_address -> servo_controllerv1_0:address
	wire         mm_interconnect_0_servo_controllerv1_0_avalon_slave_0_read;                       // mm_interconnect_0:servo_controllerv1_0_avalon_slave_0_read -> servo_controllerv1_0:read_n
	wire         mm_interconnect_0_servo_controllerv1_0_avalon_slave_0_write;                      // mm_interconnect_0:servo_controllerv1_0_avalon_slave_0_write -> servo_controllerv1_0:write_n
	wire  [31:0] mm_interconnect_0_servo_controllerv1_0_avalon_slave_0_writedata;                  // mm_interconnect_0:servo_controllerv1_0_avalon_slave_0_writedata -> servo_controllerv1_0:writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_control_slave_readdata;                              // sysid_qsys:readdata -> mm_interconnect_0:sysid_qsys_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_control_slave_address;                               // mm_interconnect_0:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire  [31:0] mm_interconnect_0_nios2_qsys_debug_mem_slave_readdata;                            // nios2_qsys:debug_mem_slave_readdata -> mm_interconnect_0:nios2_qsys_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_qsys_debug_mem_slave_waitrequest;                         // nios2_qsys:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_qsys_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_qsys_debug_mem_slave_debugaccess;                         // mm_interconnect_0:nios2_qsys_debug_mem_slave_debugaccess -> nios2_qsys:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_qsys_debug_mem_slave_address;                             // mm_interconnect_0:nios2_qsys_debug_mem_slave_address -> nios2_qsys:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_qsys_debug_mem_slave_read;                                // mm_interconnect_0:nios2_qsys_debug_mem_slave_read -> nios2_qsys:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_qsys_debug_mem_slave_byteenable;                          // mm_interconnect_0:nios2_qsys_debug_mem_slave_byteenable -> nios2_qsys:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_qsys_debug_mem_slave_write;                               // mm_interconnect_0:nios2_qsys_debug_mem_slave_write -> nios2_qsys:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_qsys_debug_mem_slave_writedata;                           // mm_interconnect_0:nios2_qsys_debug_mem_slave_writedata -> nios2_qsys:debug_mem_slave_writedata
	wire         mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_chipselect;           // mm_interconnect_0:epcs_flash_controller_0_epcs_control_port_chipselect -> epcs_flash_controller_0:chipselect
	wire  [31:0] mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_readdata;             // epcs_flash_controller_0:readdata -> mm_interconnect_0:epcs_flash_controller_0_epcs_control_port_readdata
	wire   [8:0] mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_address;              // mm_interconnect_0:epcs_flash_controller_0_epcs_control_port_address -> epcs_flash_controller_0:address
	wire         mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_read;                 // mm_interconnect_0:epcs_flash_controller_0_epcs_control_port_read -> epcs_flash_controller_0:read_n
	wire         mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_write;                // mm_interconnect_0:epcs_flash_controller_0_epcs_control_port_write -> epcs_flash_controller_0:write_n
	wire  [31:0] mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_writedata;            // mm_interconnect_0:epcs_flash_controller_0_epcs_control_port_writedata -> epcs_flash_controller_0:writedata
	wire         mm_interconnect_0_timer_s1_chipselect;                                            // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                                              // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                                               // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_write;                                                 // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                                             // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                                            // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                                              // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                                           // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                                               // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                                                  // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                                            // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                                         // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                                                 // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                                             // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_timestamp_s1_chipselect;                                        // mm_interconnect_0:timestamp_s1_chipselect -> timestamp:chipselect
	wire  [15:0] mm_interconnect_0_timestamp_s1_readdata;                                          // timestamp:readdata -> mm_interconnect_0:timestamp_s1_readdata
	wire   [3:0] mm_interconnect_0_timestamp_s1_address;                                           // mm_interconnect_0:timestamp_s1_address -> timestamp:address
	wire         mm_interconnect_0_timestamp_s1_write;                                             // mm_interconnect_0:timestamp_s1_write -> timestamp:write_n
	wire  [15:0] mm_interconnect_0_timestamp_s1_writedata;                                         // mm_interconnect_0:timestamp_s1_writedata -> timestamp:writedata
	wire  [31:0] mm_interconnect_0_uart_rs485_s1_readdata;                                         // uart_rs485:readdata -> mm_interconnect_0:uart_rs485_s1_readdata
	wire   [3:0] mm_interconnect_0_uart_rs485_s1_address;                                          // mm_interconnect_0:uart_rs485_s1_address -> uart_rs485:address
	wire         mm_interconnect_0_uart_rs485_s1_read;                                             // mm_interconnect_0:uart_rs485_s1_read -> uart_rs485:read_n
	wire         mm_interconnect_0_uart_rs485_s1_write;                                            // mm_interconnect_0:uart_rs485_s1_write -> uart_rs485:write_n
	wire  [31:0] mm_interconnect_0_uart_rs485_s1_writedata;                                        // mm_interconnect_0:uart_rs485_s1_writedata -> uart_rs485:writedata
	wire  [31:0] mm_interconnect_0_tmp101_s1_readdata;                                             // tmp101:readdata -> mm_interconnect_0:tmp101_s1_readdata
	wire   [3:0] mm_interconnect_0_tmp101_s1_address;                                              // mm_interconnect_0:tmp101_s1_address -> tmp101:address
	wire         mm_interconnect_0_tmp101_s1_read;                                                 // mm_interconnect_0:tmp101_s1_read -> tmp101:read_n
	wire         mm_interconnect_0_tmp101_s1_write;                                                // mm_interconnect_0:tmp101_s1_write -> tmp101:write_n
	wire  [31:0] mm_interconnect_0_tmp101_s1_writedata;                                            // mm_interconnect_0:tmp101_s1_writedata -> tmp101:writedata
	wire  [31:0] mm_interconnect_0_ltc2992_s1_readdata;                                            // ltc2992:readdata -> mm_interconnect_0:ltc2992_s1_readdata
	wire   [3:0] mm_interconnect_0_ltc2992_s1_address;                                             // mm_interconnect_0:ltc2992_s1_address -> ltc2992:address
	wire         mm_interconnect_0_ltc2992_s1_read;                                                // mm_interconnect_0:ltc2992_s1_read -> ltc2992:read_n
	wire         mm_interconnect_0_ltc2992_s1_write;                                               // mm_interconnect_0:ltc2992_s1_write -> ltc2992:write_n
	wire  [31:0] mm_interconnect_0_ltc2992_s1_writedata;                                           // mm_interconnect_0:ltc2992_s1_writedata -> ltc2992:writedata
	wire         mm_interconnect_0_tc_instruct_mem_s2_chipselect;                                  // mm_interconnect_0:tc_instruct_mem_s2_chipselect -> tc_instruct_mem:chipselect2
	wire  [31:0] mm_interconnect_0_tc_instruct_mem_s2_readdata;                                    // tc_instruct_mem:readdata2 -> mm_interconnect_0:tc_instruct_mem_s2_readdata
	wire  [12:0] mm_interconnect_0_tc_instruct_mem_s2_address;                                     // mm_interconnect_0:tc_instruct_mem_s2_address -> tc_instruct_mem:address2
	wire   [3:0] mm_interconnect_0_tc_instruct_mem_s2_byteenable;                                  // mm_interconnect_0:tc_instruct_mem_s2_byteenable -> tc_instruct_mem:byteenable2
	wire         mm_interconnect_0_tc_instruct_mem_s2_write;                                       // mm_interconnect_0:tc_instruct_mem_s2_write -> tc_instruct_mem:write2
	wire  [31:0] mm_interconnect_0_tc_instruct_mem_s2_writedata;                                   // mm_interconnect_0:tc_instruct_mem_s2_writedata -> tc_instruct_mem:writedata2
	wire         mm_interconnect_0_tc_instruct_mem_s2_clken;                                       // mm_interconnect_0:tc_instruct_mem_s2_clken -> tc_instruct_mem:clken2
	wire         mm_interconnect_0_boot_rom_s2_chipselect;                                         // mm_interconnect_0:boot_rom_s2_chipselect -> boot_rom:chipselect2
	wire  [31:0] mm_interconnect_0_boot_rom_s2_readdata;                                           // boot_rom:readdata2 -> mm_interconnect_0:boot_rom_s2_readdata
	wire  [10:0] mm_interconnect_0_boot_rom_s2_address;                                            // mm_interconnect_0:boot_rom_s2_address -> boot_rom:address2
	wire   [3:0] mm_interconnect_0_boot_rom_s2_byteenable;                                         // mm_interconnect_0:boot_rom_s2_byteenable -> boot_rom:byteenable2
	wire         mm_interconnect_0_boot_rom_s2_write;                                              // mm_interconnect_0:boot_rom_s2_write -> boot_rom:write2
	wire  [31:0] mm_interconnect_0_boot_rom_s2_writedata;                                          // mm_interconnect_0:boot_rom_s2_writedata -> boot_rom:writedata2
	wire         mm_interconnect_0_boot_rom_s2_clken;                                              // mm_interconnect_0:boot_rom_s2_clken -> boot_rom:clken2
	wire  [31:0] nios2_qsys_tightly_coupled_instruction_master_0_readdata;                         // mm_interconnect_1:nios2_qsys_tightly_coupled_instruction_master_0_readdata -> nios2_qsys:itcm0_readdata
	wire  [27:0] nios2_qsys_tightly_coupled_instruction_master_0_address;                          // nios2_qsys:itcm0_address -> mm_interconnect_1:nios2_qsys_tightly_coupled_instruction_master_0_address
	wire         nios2_qsys_tightly_coupled_instruction_master_0_read;                             // nios2_qsys:itcm0_read -> mm_interconnect_1:nios2_qsys_tightly_coupled_instruction_master_0_read
	wire         nios2_qsys_tightly_coupled_instruction_master_0_clken;                            // nios2_qsys:itcm0_clken -> mm_interconnect_1:nios2_qsys_tightly_coupled_instruction_master_0_clken
	wire         mm_interconnect_1_tc_instruct_mem_s1_chipselect;                                  // mm_interconnect_1:tc_instruct_mem_s1_chipselect -> tc_instruct_mem:chipselect
	wire  [31:0] mm_interconnect_1_tc_instruct_mem_s1_readdata;                                    // tc_instruct_mem:readdata -> mm_interconnect_1:tc_instruct_mem_s1_readdata
	wire  [12:0] mm_interconnect_1_tc_instruct_mem_s1_address;                                     // mm_interconnect_1:tc_instruct_mem_s1_address -> tc_instruct_mem:address
	wire   [3:0] mm_interconnect_1_tc_instruct_mem_s1_byteenable;                                  // mm_interconnect_1:tc_instruct_mem_s1_byteenable -> tc_instruct_mem:byteenable
	wire         mm_interconnect_1_tc_instruct_mem_s1_write;                                       // mm_interconnect_1:tc_instruct_mem_s1_write -> tc_instruct_mem:write
	wire  [31:0] mm_interconnect_1_tc_instruct_mem_s1_writedata;                                   // mm_interconnect_1:tc_instruct_mem_s1_writedata -> tc_instruct_mem:writedata
	wire         mm_interconnect_1_tc_instruct_mem_s1_clken;                                       // mm_interconnect_1:tc_instruct_mem_s1_clken -> tc_instruct_mem:clken
	wire  [31:0] nios2_qsys_tightly_coupled_instruction_master_1_readdata;                         // mm_interconnect_2:nios2_qsys_tightly_coupled_instruction_master_1_readdata -> nios2_qsys:itcm1_readdata
	wire  [27:0] nios2_qsys_tightly_coupled_instruction_master_1_address;                          // nios2_qsys:itcm1_address -> mm_interconnect_2:nios2_qsys_tightly_coupled_instruction_master_1_address
	wire         nios2_qsys_tightly_coupled_instruction_master_1_read;                             // nios2_qsys:itcm1_read -> mm_interconnect_2:nios2_qsys_tightly_coupled_instruction_master_1_read
	wire         nios2_qsys_tightly_coupled_instruction_master_1_clken;                            // nios2_qsys:itcm1_clken -> mm_interconnect_2:nios2_qsys_tightly_coupled_instruction_master_1_clken
	wire         mm_interconnect_2_boot_rom_s1_chipselect;                                         // mm_interconnect_2:boot_rom_s1_chipselect -> boot_rom:chipselect
	wire  [31:0] mm_interconnect_2_boot_rom_s1_readdata;                                           // boot_rom:readdata -> mm_interconnect_2:boot_rom_s1_readdata
	wire  [10:0] mm_interconnect_2_boot_rom_s1_address;                                            // mm_interconnect_2:boot_rom_s1_address -> boot_rom:address
	wire   [3:0] mm_interconnect_2_boot_rom_s1_byteenable;                                         // mm_interconnect_2:boot_rom_s1_byteenable -> boot_rom:byteenable
	wire         mm_interconnect_2_boot_rom_s1_write;                                              // mm_interconnect_2:boot_rom_s1_write -> boot_rom:write
	wire  [31:0] mm_interconnect_2_boot_rom_s1_writedata;                                          // mm_interconnect_2:boot_rom_s1_writedata -> boot_rom:writedata
	wire         mm_interconnect_2_boot_rom_s1_clken;                                              // mm_interconnect_2:boot_rom_s1_clken -> boot_rom:clken
	wire         irq_mapper_receiver0_irq;                                                         // servo_controllerv1_0:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                         // uart_rs485:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                                         // timer:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                                         // jtag_uart:av_irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                                         // epcs_flash_controller_0:irq -> irq_mapper:receiver4_irq
	wire         irq_mapper_receiver5_irq;                                                         // timestamp:irq -> irq_mapper:receiver5_irq
	wire  [31:0] nios2_qsys_irq_irq;                                                               // irq_mapper:sender_irq -> nios2_qsys:irq
	wire         rst_controller_reset_out_reset;                                                   // rst_controller:reset_out -> [boot_rom:reset, boot_rom:reset2, epcs_flash_controller_0:reset_n, jtag_uart:rst_n, mm_interconnect_0:jtag_uart_reset_reset_bridge_in_reset_reset, mm_interconnect_2:boot_rom_reset1_reset_bridge_in_reset_reset, rst_translator:in_reset, sdram:reset_n, sysid_qsys:reset_n, timer:reset_n]
	wire         rst_controller_reset_out_reset_req;                                               // rst_controller:reset_req -> [boot_rom:reset_req, boot_rom:reset_req2, epcs_flash_controller_0:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                                               // rst_controller_001:reset_out -> [irq_mapper:reset, ltc2992:reset_n, mm_interconnect_0:nios2_qsys_reset_reset_bridge_in_reset_reset, mm_interconnect_1:nios2_qsys_reset_reset_bridge_in_reset_reset, mm_interconnect_2:nios2_qsys_reset_reset_bridge_in_reset_reset, nios2_qsys:reset_n, rst_translator_001:in_reset, servo_controllerv1_0:reset_n, tc_instruct_mem:reset, tc_instruct_mem:reset2, timestamp:reset_n, tmp101:reset_n, uart_rs485:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                                           // rst_controller_001:reset_req -> [nios2_qsys:reset_req, rst_translator_001:reset_req_in, tc_instruct_mem:reset_req, tc_instruct_mem:reset_req2]
	wire         nios2_qsys_debug_reset_request_reset;                                             // nios2_qsys:debug_reset_request -> rst_controller_001:reset_in1

	DE0_CV_QSYS_boot_rom boot_rom (
		.clk         (pll_outclk0_clk),                          //   clk1.clk
		.address     (mm_interconnect_2_boot_rom_s1_address),    //     s1.address
		.clken       (mm_interconnect_2_boot_rom_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_2_boot_rom_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_2_boot_rom_s1_write),      //       .write
		.readdata    (mm_interconnect_2_boot_rom_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_2_boot_rom_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_2_boot_rom_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),           // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),       //       .reset_req
		.address2    (mm_interconnect_0_boot_rom_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_boot_rom_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_boot_rom_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_boot_rom_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_boot_rom_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_boot_rom_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_boot_rom_s2_byteenable), //       .byteenable
		.clk2        (pll_outclk0_clk),                          //   clk2.clk
		.reset2      (rst_controller_reset_out_reset),           // reset2.reset
		.reset_req2  (rst_controller_reset_out_reset_req),       //       .reset_req
		.freeze      (1'b0)                                      // (terminated)
	);

	DE0_CV_QSYS_epcs_flash_controller_0 epcs_flash_controller_0 (
		.clk        (pll_outclk0_clk),                                                        //               clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                                        //             reset.reset_n
		.reset_req  (rst_controller_reset_out_reset_req),                                     //                  .reset_req
		.address    (mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_address),    // epcs_control_port.address
		.chipselect (mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_chipselect), //                  .chipselect
		.read_n     (~mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_read),      //                  .read_n
		.readdata   (mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_readdata),   //                  .readdata
		.write_n    (~mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_write),     //                  .write_n
		.writedata  (mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_writedata),  //                  .writedata
		.irq        (irq_mapper_receiver4_irq)                                                //               irq.irq
	);

	DE0_CV_QSYS_jtag_uart jtag_uart (
		.clk            (pll_outclk0_clk),                                           //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver3_irq)                                   //               irq.irq
	);

	avl_ltc2992 #(
		.FREQ_CLK (100000000),
		.BUS_CLK  (10000)
	) ltc2992 (
		.clk       (pll_outclk0_clk),                        // clock.clk
		.reset_n   (~rst_controller_001_reset_out_reset),    // reset.reset_n
		.address   (mm_interconnect_0_ltc2992_s1_address),   //    s1.address
		.writedata (mm_interconnect_0_ltc2992_s1_writedata), //      .writedata
		.write_n   (~mm_interconnect_0_ltc2992_s1_write),    //      .write_n
		.read_n    (~mm_interconnect_0_ltc2992_s1_read),     //      .read_n
		.readdata  (mm_interconnect_0_ltc2992_s1_readdata),  //      .readdata
		.sda_t     (ltc2992_i2c_sda_t),                      //   i2c.sda_t
		.scl_t     (ltc2992_i2c_scl_t),                      //      .scl_t
		.sda_i     (ltc2992_i2c_sda_i),                      //      .sda_i
		.scl_i     (ltc2992_i2c_scl_i)                       //      .scl_i
	);

	DE0_CV_QSYS_nios2_qsys nios2_qsys (
		.clk                                 (pll_outclk0_clk),                                          //                                  clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                      //                                reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),                   //                                     .reset_req
		.d_address                           (nios2_qsys_data_master_address),                           //                          data_master.address
		.d_byteenable                        (nios2_qsys_data_master_byteenable),                        //                                     .byteenable
		.d_read                              (nios2_qsys_data_master_read),                              //                                     .read
		.d_readdata                          (nios2_qsys_data_master_readdata),                          //                                     .readdata
		.d_waitrequest                       (nios2_qsys_data_master_waitrequest),                       //                                     .waitrequest
		.d_write                             (nios2_qsys_data_master_write),                             //                                     .write
		.d_writedata                         (nios2_qsys_data_master_writedata),                         //                                     .writedata
		.d_readdatavalid                     (nios2_qsys_data_master_readdatavalid),                     //                                     .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_qsys_data_master_debugaccess),                       //                                     .debugaccess
		.i_address                           (nios2_qsys_instruction_master_address),                    //                   instruction_master.address
		.i_read                              (nios2_qsys_instruction_master_read),                       //                                     .read
		.i_readdata                          (nios2_qsys_instruction_master_readdata),                   //                                     .readdata
		.i_waitrequest                       (nios2_qsys_instruction_master_waitrequest),                //                                     .waitrequest
		.i_readdatavalid                     (nios2_qsys_instruction_master_readdatavalid),              //                                     .readdatavalid
		.itcm0_readdata                      (nios2_qsys_tightly_coupled_instruction_master_0_readdata), // tightly_coupled_instruction_master_0.readdata
		.itcm0_address                       (nios2_qsys_tightly_coupled_instruction_master_0_address),  //                                     .address
		.itcm0_read                          (nios2_qsys_tightly_coupled_instruction_master_0_read),     //                                     .read
		.itcm0_clken                         (nios2_qsys_tightly_coupled_instruction_master_0_clken),    //                                     .clken
		.itcm1_readdata                      (nios2_qsys_tightly_coupled_instruction_master_1_readdata), // tightly_coupled_instruction_master_1.readdata
		.itcm1_address                       (nios2_qsys_tightly_coupled_instruction_master_1_address),  //                                     .address
		.itcm1_read                          (nios2_qsys_tightly_coupled_instruction_master_1_read),     //                                     .read
		.itcm1_clken                         (nios2_qsys_tightly_coupled_instruction_master_1_clken),    //                                     .clken
		.irq                                 (nios2_qsys_irq_irq),                                       //                                  irq.irq
		.debug_reset_request                 (nios2_qsys_debug_reset_request_reset),                     //                  debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_qsys_debug_mem_slave_address),     //                      debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_qsys_debug_mem_slave_byteenable),  //                                     .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_qsys_debug_mem_slave_debugaccess), //                                     .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_qsys_debug_mem_slave_read),        //                                     .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_qsys_debug_mem_slave_readdata),    //                                     .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_qsys_debug_mem_slave_waitrequest), //                                     .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_qsys_debug_mem_slave_write),       //                                     .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_qsys_debug_mem_slave_writedata),   //                                     .writedata
		.A_ci_multi_done                     (nios2_qsys_custom_instruction_master_done),                //            custom_instruction_master.done
		.A_ci_multi_result                   (nios2_qsys_custom_instruction_master_multi_result),        //                                     .multi_result
		.A_ci_multi_a                        (nios2_qsys_custom_instruction_master_multi_a),             //                                     .multi_a
		.A_ci_multi_b                        (nios2_qsys_custom_instruction_master_multi_b),             //                                     .multi_b
		.A_ci_multi_c                        (nios2_qsys_custom_instruction_master_multi_c),             //                                     .multi_c
		.A_ci_multi_clk_en                   (nios2_qsys_custom_instruction_master_clk_en),              //                                     .clk_en
		.A_ci_multi_clock                    (nios2_qsys_custom_instruction_master_clk),                 //                                     .clk
		.A_ci_multi_reset                    (nios2_qsys_custom_instruction_master_reset),               //                                     .reset
		.A_ci_multi_reset_req                (nios2_qsys_custom_instruction_master_reset_req),           //                                     .reset_req
		.A_ci_multi_dataa                    (nios2_qsys_custom_instruction_master_multi_dataa),         //                                     .multi_dataa
		.A_ci_multi_datab                    (nios2_qsys_custom_instruction_master_multi_datab),         //                                     .multi_datab
		.A_ci_multi_n                        (nios2_qsys_custom_instruction_master_multi_n),             //                                     .multi_n
		.A_ci_multi_readra                   (nios2_qsys_custom_instruction_master_multi_readra),        //                                     .multi_readra
		.A_ci_multi_readrb                   (nios2_qsys_custom_instruction_master_multi_readrb),        //                                     .multi_readrb
		.A_ci_multi_start                    (nios2_qsys_custom_instruction_master_start),               //                                     .start
		.A_ci_multi_writerc                  (nios2_qsys_custom_instruction_master_multi_writerc),       //                                     .multi_writerc
		.E_ci_combo_result                   (nios2_qsys_custom_instruction_master_result),              //                                     .result
		.E_ci_combo_a                        (nios2_qsys_custom_instruction_master_a),                   //                                     .a
		.E_ci_combo_b                        (nios2_qsys_custom_instruction_master_b),                   //                                     .b
		.E_ci_combo_c                        (nios2_qsys_custom_instruction_master_c),                   //                                     .c
		.E_ci_combo_dataa                    (nios2_qsys_custom_instruction_master_dataa),               //                                     .dataa
		.E_ci_combo_datab                    (nios2_qsys_custom_instruction_master_datab),               //                                     .datab
		.E_ci_combo_estatus                  (nios2_qsys_custom_instruction_master_estatus),             //                                     .estatus
		.E_ci_combo_ipending                 (nios2_qsys_custom_instruction_master_ipending),            //                                     .ipending
		.E_ci_combo_n                        (nios2_qsys_custom_instruction_master_n),                   //                                     .n
		.E_ci_combo_readra                   (nios2_qsys_custom_instruction_master_readra),              //                                     .readra
		.E_ci_combo_readrb                   (nios2_qsys_custom_instruction_master_readrb),              //                                     .readrb
		.E_ci_combo_writerc                  (nios2_qsys_custom_instruction_master_writerc)              //                                     .writerc
	);

	DE0_CV_QSYS_nios_custom_instr_floating_point_2_0 #(
		.arithmetic_present (1),
		.root_present       (1),
		.conversion_present (1),
		.comparison_present (1)
	) nios_custom_instr_floating_point_2_0 (
		.s1_dataa     (nios2_qsys_custom_instruction_master_comb_slave_translator0_ci_master_dataa),      // s1.dataa
		.s1_datab     (nios2_qsys_custom_instruction_master_comb_slave_translator0_ci_master_datab),      //   .datab
		.s1_n         (nios2_qsys_custom_instruction_master_comb_slave_translator0_ci_master_n),          //   .n
		.s1_result    (nios2_qsys_custom_instruction_master_comb_slave_translator0_ci_master_result),     //   .result
		.s2_clk       (nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_clk),       // s2.clk
		.s2_clk_en    (nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_clk_en),    //   .clk_en
		.s2_dataa     (nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_dataa),     //   .dataa
		.s2_datab     (nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_datab),     //   .datab
		.s2_n         (nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_n),         //   .n
		.s2_reset     (nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_reset),     //   .reset
		.s2_reset_req (nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_reset_req), //   .reset_req
		.s2_start     (nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_start),     //   .start
		.s2_done      (nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_done),      //   .done
		.s2_result    (nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_result)     //   .result
	);

	DE0_CV_QSYS_pll pll (
		.refclk   (clk_clk),           //  refclk.clk
		.rst      (~reset_reset_n),    //   reset.reset
		.outclk_0 (pll_outclk0_clk),   // outclk0.clk
		.outclk_1 (clk_sdram_clk),     // outclk1.clk
		.outclk_2 (clk_5m_clk),        // outclk2.clk
		.locked   (pll_locked_export)  //  locked.export
	);

	DE0_CV_QSYS_sdram sdram (
		.clk            (pll_outclk0_clk),                          //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	servo_controllerv1 #(
		.FREQ_CLK      (100000000),
		.SPI_SPEED     (1000000),
		.PWM_BASE_FREQ (10000000),
		.PWM_FREQ      (1000),
		.C_MODE0       (0),
		.C_MODE1       (0),
		.C_MODE2       (0),
		.C_MODE3       (0)
	) servo_controllerv1_0 (
		.clk        (pll_outclk0_clk),                                                 //            clock.clk
		.reset_n    (~rst_controller_001_reset_out_reset),                             //            reset.reset_n
		.address    (mm_interconnect_0_servo_controllerv1_0_avalon_slave_0_address),   //   avalon_slave_0.address
		.writedata  (mm_interconnect_0_servo_controllerv1_0_avalon_slave_0_writedata), //                 .writedata
		.write_n    (~mm_interconnect_0_servo_controllerv1_0_avalon_slave_0_write),    //                 .write_n
		.read_n     (~mm_interconnect_0_servo_controllerv1_0_avalon_slave_0_read),     //                 .read_n
		.readdata   (mm_interconnect_0_servo_controllerv1_0_avalon_slave_0_readdata),  //                 .readdata
		.spi_sclk   (servo_controllerv1_0_conduit_end_spi_sclk),                       //      conduit_end.spi_sclk
		.spi_cs     (servo_controllerv1_0_conduit_end_spi_cs),                         //                 .spi_cs
		.spi_miso   (servo_controllerv1_0_conduit_end_spi_miso),                       //                 .spi_miso
		.spi_mosi   (servo_controllerv1_0_conduit_end_spi_mosi),                       //                 .spi_mosi
		.hall_0     (servo_controllerv1_0_conduit_end_hall_0),                         //                 .hall_0
		.hall_1     (servo_controllerv1_0_conduit_end_hall_1),                         //                 .hall_1
		.hall_2     (servo_controllerv1_0_conduit_end_hall_2),                         //                 .hall_2
		.hall_3     (servo_controllerv1_0_conduit_end_hall_3),                         //                 .hall_3
		.phase_0    (servo_controllerv1_0_conduit_end_phase_0),                        //                 .phase_0
		.phase_1    (servo_controllerv1_0_conduit_end_phase_1),                        //                 .phase_1
		.phase_2    (servo_controllerv1_0_conduit_end_phase_2),                        //                 .phase_2
		.phase_3    (servo_controllerv1_0_conduit_end_phase_3),                        //                 .phase_3
		.nFault     (servo_controllerv1_0_conduit_end_nFault),                         //                 .nFault
		.drv8320_en (servo_controllerv1_0_conduit_end_drv8320_en),                     //                 .drv8320_en
		.irq        (irq_mapper_receiver0_irq)                                         // interrupt_sender.irq
	);

	DE0_CV_QSYS_sysid_qsys sysid_qsys (
		.clock    (pll_outclk0_clk),                                     //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                     //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_control_slave_address)   //              .address
	);

	DE0_CV_QSYS_tc_instruct_mem tc_instruct_mem (
		.clk         (pll_outclk0_clk),                                 //   clk1.clk
		.address     (mm_interconnect_1_tc_instruct_mem_s1_address),    //     s1.address
		.clken       (mm_interconnect_1_tc_instruct_mem_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_1_tc_instruct_mem_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_1_tc_instruct_mem_s1_write),      //       .write
		.readdata    (mm_interconnect_1_tc_instruct_mem_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_1_tc_instruct_mem_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_1_tc_instruct_mem_s1_byteenable), //       .byteenable
		.reset       (rst_controller_001_reset_out_reset),              // reset1.reset
		.reset_req   (rst_controller_001_reset_out_reset_req),          //       .reset_req
		.address2    (mm_interconnect_0_tc_instruct_mem_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_tc_instruct_mem_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_tc_instruct_mem_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_tc_instruct_mem_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_tc_instruct_mem_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_tc_instruct_mem_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_tc_instruct_mem_s2_byteenable), //       .byteenable
		.clk2        (pll_outclk0_clk),                                 //   clk2.clk
		.reset2      (rst_controller_001_reset_out_reset),              // reset2.reset
		.reset_req2  (rst_controller_001_reset_out_reset_req),          //       .reset_req
		.freeze      (1'b0)                                             // (terminated)
	);

	DE0_CV_QSYS_timer timer (
		.clk        (pll_outclk0_clk),                       //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)               //   irq.irq
	);

	DE0_CV_QSYS_timestamp timestamp (
		.clk        (pll_outclk0_clk),                           //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timestamp_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timestamp_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timestamp_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timestamp_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timestamp_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver5_irq)                   //   irq.irq
	);

	avl_tmp101 #(
		.FREQ_CLK    (100000000),
		.BUS_CLK     (100000),
		.UPDATE_FREQ (2),
		.I2C_ADDR    (0)
	) tmp101 (
		.clk       (pll_outclk0_clk),                       // clock.clk
		.reset_n   (~rst_controller_001_reset_out_reset),   // reset.reset_n
		.address   (mm_interconnect_0_tmp101_s1_address),   //    s1.address
		.writedata (mm_interconnect_0_tmp101_s1_writedata), //      .writedata
		.write_n   (~mm_interconnect_0_tmp101_s1_write),    //      .write_n
		.read_n    (~mm_interconnect_0_tmp101_s1_read),     //      .read_n
		.readdata  (mm_interconnect_0_tmp101_s1_readdata),  //      .readdata
		.sda_t     (tmp101_i2c_sda_t),                      //   i2c.sda_t
		.scl_t     (tmp101_i2c_scl_t),                      //      .scl_t
		.sda_i     (tmp101_i2c_sda_i),                      //      .sda_i
		.scl_i     (tmp101_i2c_scl_i)                       //      .scl_i
	);

	avl_fifo_uart #(
		.FREQ_CLK          (100000000),
		.BAUDRATE          (921600),
		.DATA_BIT          (8),
		.PARITY_BIT        (0),
		.STOP_BIT          (0),
		.C_RX_THRESHOLD    (32),
		.RX_FIFO_DEPTH     (7),
		.TX_FIFO_DEPTH     (12),
		.OVERSAMPLING_RATE (4),
		.RX_TIMEOUT_WORD   (4)
	) uart_rs485 (
		.clk          (pll_outclk0_clk),                           //            clock.clk
		.reset_n      (~rst_controller_001_reset_out_reset),       //            reset.reset_n
		.address      (mm_interconnect_0_uart_rs485_s1_address),   //               s1.address
		.writedata    (mm_interconnect_0_uart_rs485_s1_writedata), //                 .writedata
		.write_n      (~mm_interconnect_0_uart_rs485_s1_write),    //                 .write_n
		.read_n       (~mm_interconnect_0_uart_rs485_s1_read),     //                 .read_n
		.readdata     (mm_interconnect_0_uart_rs485_s1_readdata),  //                 .readdata
		.rxd          (uart_rs485_conduit_end_rxd),                //      conduit_end.rxd
		.txd          (uart_rs485_conduit_end_txd),                //                 .txd
		.dbg_os_pulse (uart_rs485_conduit_end_dbg_os_pulse),       //                 .dbg_os_pulse
		.irq          (irq_mapper_receiver1_irq)                   // interrupt_sender.irq
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (0)
	) nios2_qsys_custom_instruction_master_translator (
		.ci_slave_dataa            (nios2_qsys_custom_instruction_master_dataa),                                //        ci_slave.dataa
		.ci_slave_datab            (nios2_qsys_custom_instruction_master_datab),                                //                .datab
		.ci_slave_result           (nios2_qsys_custom_instruction_master_result),                               //                .result
		.ci_slave_n                (nios2_qsys_custom_instruction_master_n),                                    //                .n
		.ci_slave_readra           (nios2_qsys_custom_instruction_master_readra),                               //                .readra
		.ci_slave_readrb           (nios2_qsys_custom_instruction_master_readrb),                               //                .readrb
		.ci_slave_writerc          (nios2_qsys_custom_instruction_master_writerc),                              //                .writerc
		.ci_slave_a                (nios2_qsys_custom_instruction_master_a),                                    //                .a
		.ci_slave_b                (nios2_qsys_custom_instruction_master_b),                                    //                .b
		.ci_slave_c                (nios2_qsys_custom_instruction_master_c),                                    //                .c
		.ci_slave_ipending         (nios2_qsys_custom_instruction_master_ipending),                             //                .ipending
		.ci_slave_estatus          (nios2_qsys_custom_instruction_master_estatus),                              //                .estatus
		.ci_slave_multi_clk        (nios2_qsys_custom_instruction_master_clk),                                  //                .clk
		.ci_slave_multi_reset      (nios2_qsys_custom_instruction_master_reset),                                //                .reset
		.ci_slave_multi_clken      (nios2_qsys_custom_instruction_master_clk_en),                               //                .clk_en
		.ci_slave_multi_reset_req  (nios2_qsys_custom_instruction_master_reset_req),                            //                .reset_req
		.ci_slave_multi_start      (nios2_qsys_custom_instruction_master_start),                                //                .start
		.ci_slave_multi_done       (nios2_qsys_custom_instruction_master_done),                                 //                .done
		.ci_slave_multi_dataa      (nios2_qsys_custom_instruction_master_multi_dataa),                          //                .multi_dataa
		.ci_slave_multi_datab      (nios2_qsys_custom_instruction_master_multi_datab),                          //                .multi_datab
		.ci_slave_multi_result     (nios2_qsys_custom_instruction_master_multi_result),                         //                .multi_result
		.ci_slave_multi_n          (nios2_qsys_custom_instruction_master_multi_n),                              //                .multi_n
		.ci_slave_multi_readra     (nios2_qsys_custom_instruction_master_multi_readra),                         //                .multi_readra
		.ci_slave_multi_readrb     (nios2_qsys_custom_instruction_master_multi_readrb),                         //                .multi_readrb
		.ci_slave_multi_writerc    (nios2_qsys_custom_instruction_master_multi_writerc),                        //                .multi_writerc
		.ci_slave_multi_a          (nios2_qsys_custom_instruction_master_multi_a),                              //                .multi_a
		.ci_slave_multi_b          (nios2_qsys_custom_instruction_master_multi_b),                              //                .multi_b
		.ci_slave_multi_c          (nios2_qsys_custom_instruction_master_multi_c),                              //                .multi_c
		.comb_ci_master_dataa      (nios2_qsys_custom_instruction_master_translator_comb_ci_master_dataa),      //  comb_ci_master.dataa
		.comb_ci_master_datab      (nios2_qsys_custom_instruction_master_translator_comb_ci_master_datab),      //                .datab
		.comb_ci_master_result     (nios2_qsys_custom_instruction_master_translator_comb_ci_master_result),     //                .result
		.comb_ci_master_n          (nios2_qsys_custom_instruction_master_translator_comb_ci_master_n),          //                .n
		.comb_ci_master_readra     (nios2_qsys_custom_instruction_master_translator_comb_ci_master_readra),     //                .readra
		.comb_ci_master_readrb     (nios2_qsys_custom_instruction_master_translator_comb_ci_master_readrb),     //                .readrb
		.comb_ci_master_writerc    (nios2_qsys_custom_instruction_master_translator_comb_ci_master_writerc),    //                .writerc
		.comb_ci_master_a          (nios2_qsys_custom_instruction_master_translator_comb_ci_master_a),          //                .a
		.comb_ci_master_b          (nios2_qsys_custom_instruction_master_translator_comb_ci_master_b),          //                .b
		.comb_ci_master_c          (nios2_qsys_custom_instruction_master_translator_comb_ci_master_c),          //                .c
		.comb_ci_master_ipending   (nios2_qsys_custom_instruction_master_translator_comb_ci_master_ipending),   //                .ipending
		.comb_ci_master_estatus    (nios2_qsys_custom_instruction_master_translator_comb_ci_master_estatus),    //                .estatus
		.multi_ci_master_clk       (nios2_qsys_custom_instruction_master_translator_multi_ci_master_clk),       // multi_ci_master.clk
		.multi_ci_master_reset     (nios2_qsys_custom_instruction_master_translator_multi_ci_master_reset),     //                .reset
		.multi_ci_master_clken     (nios2_qsys_custom_instruction_master_translator_multi_ci_master_clk_en),    //                .clk_en
		.multi_ci_master_reset_req (nios2_qsys_custom_instruction_master_translator_multi_ci_master_reset_req), //                .reset_req
		.multi_ci_master_start     (nios2_qsys_custom_instruction_master_translator_multi_ci_master_start),     //                .start
		.multi_ci_master_done      (nios2_qsys_custom_instruction_master_translator_multi_ci_master_done),      //                .done
		.multi_ci_master_dataa     (nios2_qsys_custom_instruction_master_translator_multi_ci_master_dataa),     //                .dataa
		.multi_ci_master_datab     (nios2_qsys_custom_instruction_master_translator_multi_ci_master_datab),     //                .datab
		.multi_ci_master_result    (nios2_qsys_custom_instruction_master_translator_multi_ci_master_result),    //                .result
		.multi_ci_master_n         (nios2_qsys_custom_instruction_master_translator_multi_ci_master_n),         //                .n
		.multi_ci_master_readra    (nios2_qsys_custom_instruction_master_translator_multi_ci_master_readra),    //                .readra
		.multi_ci_master_readrb    (nios2_qsys_custom_instruction_master_translator_multi_ci_master_readrb),    //                .readrb
		.multi_ci_master_writerc   (nios2_qsys_custom_instruction_master_translator_multi_ci_master_writerc),   //                .writerc
		.multi_ci_master_a         (nios2_qsys_custom_instruction_master_translator_multi_ci_master_a),         //                .a
		.multi_ci_master_b         (nios2_qsys_custom_instruction_master_translator_multi_ci_master_b),         //                .b
		.multi_ci_master_c         (nios2_qsys_custom_instruction_master_translator_multi_ci_master_c)          //                .c
	);

	DE0_CV_QSYS_nios2_qsys_custom_instruction_master_comb_xconnect nios2_qsys_custom_instruction_master_comb_xconnect (
		.ci_slave_dataa      (nios2_qsys_custom_instruction_master_translator_comb_ci_master_dataa),    //   ci_slave.dataa
		.ci_slave_datab      (nios2_qsys_custom_instruction_master_translator_comb_ci_master_datab),    //           .datab
		.ci_slave_result     (nios2_qsys_custom_instruction_master_translator_comb_ci_master_result),   //           .result
		.ci_slave_n          (nios2_qsys_custom_instruction_master_translator_comb_ci_master_n),        //           .n
		.ci_slave_readra     (nios2_qsys_custom_instruction_master_translator_comb_ci_master_readra),   //           .readra
		.ci_slave_readrb     (nios2_qsys_custom_instruction_master_translator_comb_ci_master_readrb),   //           .readrb
		.ci_slave_writerc    (nios2_qsys_custom_instruction_master_translator_comb_ci_master_writerc),  //           .writerc
		.ci_slave_a          (nios2_qsys_custom_instruction_master_translator_comb_ci_master_a),        //           .a
		.ci_slave_b          (nios2_qsys_custom_instruction_master_translator_comb_ci_master_b),        //           .b
		.ci_slave_c          (nios2_qsys_custom_instruction_master_translator_comb_ci_master_c),        //           .c
		.ci_slave_ipending   (nios2_qsys_custom_instruction_master_translator_comb_ci_master_ipending), //           .ipending
		.ci_slave_estatus    (nios2_qsys_custom_instruction_master_translator_comb_ci_master_estatus),  //           .estatus
		.ci_master0_dataa    (nios2_qsys_custom_instruction_master_comb_xconnect_ci_master0_dataa),     // ci_master0.dataa
		.ci_master0_datab    (nios2_qsys_custom_instruction_master_comb_xconnect_ci_master0_datab),     //           .datab
		.ci_master0_result   (nios2_qsys_custom_instruction_master_comb_xconnect_ci_master0_result),    //           .result
		.ci_master0_n        (nios2_qsys_custom_instruction_master_comb_xconnect_ci_master0_n),         //           .n
		.ci_master0_readra   (nios2_qsys_custom_instruction_master_comb_xconnect_ci_master0_readra),    //           .readra
		.ci_master0_readrb   (nios2_qsys_custom_instruction_master_comb_xconnect_ci_master0_readrb),    //           .readrb
		.ci_master0_writerc  (nios2_qsys_custom_instruction_master_comb_xconnect_ci_master0_writerc),   //           .writerc
		.ci_master0_a        (nios2_qsys_custom_instruction_master_comb_xconnect_ci_master0_a),         //           .a
		.ci_master0_b        (nios2_qsys_custom_instruction_master_comb_xconnect_ci_master0_b),         //           .b
		.ci_master0_c        (nios2_qsys_custom_instruction_master_comb_xconnect_ci_master0_c),         //           .c
		.ci_master0_ipending (nios2_qsys_custom_instruction_master_comb_xconnect_ci_master0_ipending),  //           .ipending
		.ci_master0_estatus  (nios2_qsys_custom_instruction_master_comb_xconnect_ci_master0_estatus)    //           .estatus
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (4),
		.USE_DONE         (0),
		.NUM_FIXED_CYCLES (0)
	) nios2_qsys_custom_instruction_master_comb_slave_translator0 (
		.ci_slave_dataa      (nios2_qsys_custom_instruction_master_comb_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (nios2_qsys_custom_instruction_master_comb_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (nios2_qsys_custom_instruction_master_comb_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (nios2_qsys_custom_instruction_master_comb_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (nios2_qsys_custom_instruction_master_comb_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (nios2_qsys_custom_instruction_master_comb_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (nios2_qsys_custom_instruction_master_comb_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (nios2_qsys_custom_instruction_master_comb_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (nios2_qsys_custom_instruction_master_comb_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (nios2_qsys_custom_instruction_master_comb_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (nios2_qsys_custom_instruction_master_comb_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (nios2_qsys_custom_instruction_master_comb_xconnect_ci_master0_estatus),        //          .estatus
		.ci_master_dataa     (nios2_qsys_custom_instruction_master_comb_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (nios2_qsys_custom_instruction_master_comb_slave_translator0_ci_master_datab),  //          .datab
		.ci_master_result    (nios2_qsys_custom_instruction_master_comb_slave_translator0_ci_master_result), //          .result
		.ci_master_n         (nios2_qsys_custom_instruction_master_comb_slave_translator0_ci_master_n),      //          .n
		.ci_master_readra    (),                                                                             // (terminated)
		.ci_master_readrb    (),                                                                             // (terminated)
		.ci_master_writerc   (),                                                                             // (terminated)
		.ci_master_a         (),                                                                             // (terminated)
		.ci_master_b         (),                                                                             // (terminated)
		.ci_master_c         (),                                                                             // (terminated)
		.ci_master_ipending  (),                                                                             // (terminated)
		.ci_master_estatus   (),                                                                             // (terminated)
		.ci_master_clk       (),                                                                             // (terminated)
		.ci_master_clken     (),                                                                             // (terminated)
		.ci_master_reset_req (),                                                                             // (terminated)
		.ci_master_reset     (),                                                                             // (terminated)
		.ci_master_start     (),                                                                             // (terminated)
		.ci_master_done      (1'b0),                                                                         // (terminated)
		.ci_slave_clk        (1'b0),                                                                         // (terminated)
		.ci_slave_clken      (1'b0),                                                                         // (terminated)
		.ci_slave_reset_req  (1'b0),                                                                         // (terminated)
		.ci_slave_reset      (1'b0),                                                                         // (terminated)
		.ci_slave_start      (1'b0),                                                                         // (terminated)
		.ci_slave_done       ()                                                                              // (terminated)
	);

	DE0_CV_QSYS_nios2_qsys_custom_instruction_master_multi_xconnect nios2_qsys_custom_instruction_master_multi_xconnect (
		.ci_slave_dataa       (nios2_qsys_custom_instruction_master_translator_multi_ci_master_dataa),     //   ci_slave.dataa
		.ci_slave_datab       (nios2_qsys_custom_instruction_master_translator_multi_ci_master_datab),     //           .datab
		.ci_slave_result      (nios2_qsys_custom_instruction_master_translator_multi_ci_master_result),    //           .result
		.ci_slave_n           (nios2_qsys_custom_instruction_master_translator_multi_ci_master_n),         //           .n
		.ci_slave_readra      (nios2_qsys_custom_instruction_master_translator_multi_ci_master_readra),    //           .readra
		.ci_slave_readrb      (nios2_qsys_custom_instruction_master_translator_multi_ci_master_readrb),    //           .readrb
		.ci_slave_writerc     (nios2_qsys_custom_instruction_master_translator_multi_ci_master_writerc),   //           .writerc
		.ci_slave_a           (nios2_qsys_custom_instruction_master_translator_multi_ci_master_a),         //           .a
		.ci_slave_b           (nios2_qsys_custom_instruction_master_translator_multi_ci_master_b),         //           .b
		.ci_slave_c           (nios2_qsys_custom_instruction_master_translator_multi_ci_master_c),         //           .c
		.ci_slave_ipending    (),                                                                          //           .ipending
		.ci_slave_estatus     (),                                                                          //           .estatus
		.ci_slave_clk         (nios2_qsys_custom_instruction_master_translator_multi_ci_master_clk),       //           .clk
		.ci_slave_reset       (nios2_qsys_custom_instruction_master_translator_multi_ci_master_reset),     //           .reset
		.ci_slave_clken       (nios2_qsys_custom_instruction_master_translator_multi_ci_master_clk_en),    //           .clk_en
		.ci_slave_reset_req   (nios2_qsys_custom_instruction_master_translator_multi_ci_master_reset_req), //           .reset_req
		.ci_slave_start       (nios2_qsys_custom_instruction_master_translator_multi_ci_master_start),     //           .start
		.ci_slave_done        (nios2_qsys_custom_instruction_master_translator_multi_ci_master_done),      //           .done
		.ci_master0_dataa     (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_dataa),      // ci_master0.dataa
		.ci_master0_datab     (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_datab),      //           .datab
		.ci_master0_result    (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_result),     //           .result
		.ci_master0_n         (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_n),          //           .n
		.ci_master0_readra    (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_readra),     //           .readra
		.ci_master0_readrb    (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_readrb),     //           .readrb
		.ci_master0_writerc   (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_writerc),    //           .writerc
		.ci_master0_a         (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_a),          //           .a
		.ci_master0_b         (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_b),          //           .b
		.ci_master0_c         (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_c),          //           .c
		.ci_master0_ipending  (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_ipending),   //           .ipending
		.ci_master0_estatus   (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_estatus),    //           .estatus
		.ci_master0_clk       (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_clk),        //           .clk
		.ci_master0_reset     (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_reset),      //           .reset
		.ci_master0_clken     (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_clk_en),     //           .clk_en
		.ci_master0_reset_req (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_reset_req),  //           .reset_req
		.ci_master0_start     (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_start),      //           .start
		.ci_master0_done      (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_done)        //           .done
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (3),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (1)
	) nios2_qsys_custom_instruction_master_multi_slave_translator0 (
		.ci_slave_dataa      (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_dataa),             //  ci_slave.dataa
		.ci_slave_datab      (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_datab),             //          .datab
		.ci_slave_result     (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_result),            //          .result
		.ci_slave_n          (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_n),                 //          .n
		.ci_slave_readra     (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_readra),            //          .readra
		.ci_slave_readrb     (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_readrb),            //          .readrb
		.ci_slave_writerc    (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_writerc),           //          .writerc
		.ci_slave_a          (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_a),                 //          .a
		.ci_slave_b          (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_b),                 //          .b
		.ci_slave_c          (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_c),                 //          .c
		.ci_slave_ipending   (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_ipending),          //          .ipending
		.ci_slave_estatus    (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_estatus),           //          .estatus
		.ci_slave_clk        (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_clk),               //          .clk
		.ci_slave_clken      (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_clk_en),            //          .clk_en
		.ci_slave_reset_req  (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_reset_req),         //          .reset_req
		.ci_slave_reset      (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_reset),             //          .reset
		.ci_slave_start      (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_start),             //          .start
		.ci_slave_done       (nios2_qsys_custom_instruction_master_multi_xconnect_ci_master0_done),              //          .done
		.ci_master_dataa     (nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_dataa),     // ci_master.dataa
		.ci_master_datab     (nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_datab),     //          .datab
		.ci_master_result    (nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_result),    //          .result
		.ci_master_n         (nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_n),         //          .n
		.ci_master_clk       (nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_clk),       //          .clk
		.ci_master_clken     (nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_clk_en),    //          .clk_en
		.ci_master_reset_req (nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_reset_req), //          .reset_req
		.ci_master_reset     (nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_reset),     //          .reset
		.ci_master_start     (nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_start),     //          .start
		.ci_master_done      (nios2_qsys_custom_instruction_master_multi_slave_translator0_ci_master_done),      //          .done
		.ci_master_readra    (),                                                                                 // (terminated)
		.ci_master_readrb    (),                                                                                 // (terminated)
		.ci_master_writerc   (),                                                                                 // (terminated)
		.ci_master_a         (),                                                                                 // (terminated)
		.ci_master_b         (),                                                                                 // (terminated)
		.ci_master_c         (),                                                                                 // (terminated)
		.ci_master_ipending  (),                                                                                 // (terminated)
		.ci_master_estatus   ()                                                                                  // (terminated)
	);

	DE0_CV_QSYS_mm_interconnect_0 mm_interconnect_0 (
		.pll_outclk0_clk                                      (pll_outclk0_clk),                                                        //                               pll_outclk0.clk
		.jtag_uart_reset_reset_bridge_in_reset_reset          (rst_controller_reset_out_reset),                                         //     jtag_uart_reset_reset_bridge_in_reset.reset
		.nios2_qsys_reset_reset_bridge_in_reset_reset         (rst_controller_001_reset_out_reset),                                     //    nios2_qsys_reset_reset_bridge_in_reset.reset
		.nios2_qsys_data_master_address                       (nios2_qsys_data_master_address),                                         //                    nios2_qsys_data_master.address
		.nios2_qsys_data_master_waitrequest                   (nios2_qsys_data_master_waitrequest),                                     //                                          .waitrequest
		.nios2_qsys_data_master_byteenable                    (nios2_qsys_data_master_byteenable),                                      //                                          .byteenable
		.nios2_qsys_data_master_read                          (nios2_qsys_data_master_read),                                            //                                          .read
		.nios2_qsys_data_master_readdata                      (nios2_qsys_data_master_readdata),                                        //                                          .readdata
		.nios2_qsys_data_master_readdatavalid                 (nios2_qsys_data_master_readdatavalid),                                   //                                          .readdatavalid
		.nios2_qsys_data_master_write                         (nios2_qsys_data_master_write),                                           //                                          .write
		.nios2_qsys_data_master_writedata                     (nios2_qsys_data_master_writedata),                                       //                                          .writedata
		.nios2_qsys_data_master_debugaccess                   (nios2_qsys_data_master_debugaccess),                                     //                                          .debugaccess
		.nios2_qsys_instruction_master_address                (nios2_qsys_instruction_master_address),                                  //             nios2_qsys_instruction_master.address
		.nios2_qsys_instruction_master_waitrequest            (nios2_qsys_instruction_master_waitrequest),                              //                                          .waitrequest
		.nios2_qsys_instruction_master_read                   (nios2_qsys_instruction_master_read),                                     //                                          .read
		.nios2_qsys_instruction_master_readdata               (nios2_qsys_instruction_master_readdata),                                 //                                          .readdata
		.nios2_qsys_instruction_master_readdatavalid          (nios2_qsys_instruction_master_readdatavalid),                            //                                          .readdatavalid
		.boot_rom_s2_address                                  (mm_interconnect_0_boot_rom_s2_address),                                  //                               boot_rom_s2.address
		.boot_rom_s2_write                                    (mm_interconnect_0_boot_rom_s2_write),                                    //                                          .write
		.boot_rom_s2_readdata                                 (mm_interconnect_0_boot_rom_s2_readdata),                                 //                                          .readdata
		.boot_rom_s2_writedata                                (mm_interconnect_0_boot_rom_s2_writedata),                                //                                          .writedata
		.boot_rom_s2_byteenable                               (mm_interconnect_0_boot_rom_s2_byteenable),                               //                                          .byteenable
		.boot_rom_s2_chipselect                               (mm_interconnect_0_boot_rom_s2_chipselect),                               //                                          .chipselect
		.boot_rom_s2_clken                                    (mm_interconnect_0_boot_rom_s2_clken),                                    //                                          .clken
		.epcs_flash_controller_0_epcs_control_port_address    (mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_address),    // epcs_flash_controller_0_epcs_control_port.address
		.epcs_flash_controller_0_epcs_control_port_write      (mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_write),      //                                          .write
		.epcs_flash_controller_0_epcs_control_port_read       (mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_read),       //                                          .read
		.epcs_flash_controller_0_epcs_control_port_readdata   (mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_readdata),   //                                          .readdata
		.epcs_flash_controller_0_epcs_control_port_writedata  (mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_writedata),  //                                          .writedata
		.epcs_flash_controller_0_epcs_control_port_chipselect (mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_chipselect), //                                          .chipselect
		.jtag_uart_avalon_jtag_slave_address                  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),                  //               jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),                    //                                          .write
		.jtag_uart_avalon_jtag_slave_read                     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),                     //                                          .read
		.jtag_uart_avalon_jtag_slave_readdata                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),                 //                                          .readdata
		.jtag_uart_avalon_jtag_slave_writedata                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),                //                                          .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),              //                                          .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),               //                                          .chipselect
		.ltc2992_s1_address                                   (mm_interconnect_0_ltc2992_s1_address),                                   //                                ltc2992_s1.address
		.ltc2992_s1_write                                     (mm_interconnect_0_ltc2992_s1_write),                                     //                                          .write
		.ltc2992_s1_read                                      (mm_interconnect_0_ltc2992_s1_read),                                      //                                          .read
		.ltc2992_s1_readdata                                  (mm_interconnect_0_ltc2992_s1_readdata),                                  //                                          .readdata
		.ltc2992_s1_writedata                                 (mm_interconnect_0_ltc2992_s1_writedata),                                 //                                          .writedata
		.nios2_qsys_debug_mem_slave_address                   (mm_interconnect_0_nios2_qsys_debug_mem_slave_address),                   //                nios2_qsys_debug_mem_slave.address
		.nios2_qsys_debug_mem_slave_write                     (mm_interconnect_0_nios2_qsys_debug_mem_slave_write),                     //                                          .write
		.nios2_qsys_debug_mem_slave_read                      (mm_interconnect_0_nios2_qsys_debug_mem_slave_read),                      //                                          .read
		.nios2_qsys_debug_mem_slave_readdata                  (mm_interconnect_0_nios2_qsys_debug_mem_slave_readdata),                  //                                          .readdata
		.nios2_qsys_debug_mem_slave_writedata                 (mm_interconnect_0_nios2_qsys_debug_mem_slave_writedata),                 //                                          .writedata
		.nios2_qsys_debug_mem_slave_byteenable                (mm_interconnect_0_nios2_qsys_debug_mem_slave_byteenable),                //                                          .byteenable
		.nios2_qsys_debug_mem_slave_waitrequest               (mm_interconnect_0_nios2_qsys_debug_mem_slave_waitrequest),               //                                          .waitrequest
		.nios2_qsys_debug_mem_slave_debugaccess               (mm_interconnect_0_nios2_qsys_debug_mem_slave_debugaccess),               //                                          .debugaccess
		.sdram_s1_address                                     (mm_interconnect_0_sdram_s1_address),                                     //                                  sdram_s1.address
		.sdram_s1_write                                       (mm_interconnect_0_sdram_s1_write),                                       //                                          .write
		.sdram_s1_read                                        (mm_interconnect_0_sdram_s1_read),                                        //                                          .read
		.sdram_s1_readdata                                    (mm_interconnect_0_sdram_s1_readdata),                                    //                                          .readdata
		.sdram_s1_writedata                                   (mm_interconnect_0_sdram_s1_writedata),                                   //                                          .writedata
		.sdram_s1_byteenable                                  (mm_interconnect_0_sdram_s1_byteenable),                                  //                                          .byteenable
		.sdram_s1_readdatavalid                               (mm_interconnect_0_sdram_s1_readdatavalid),                               //                                          .readdatavalid
		.sdram_s1_waitrequest                                 (mm_interconnect_0_sdram_s1_waitrequest),                                 //                                          .waitrequest
		.sdram_s1_chipselect                                  (mm_interconnect_0_sdram_s1_chipselect),                                  //                                          .chipselect
		.servo_controllerv1_0_avalon_slave_0_address          (mm_interconnect_0_servo_controllerv1_0_avalon_slave_0_address),          //       servo_controllerv1_0_avalon_slave_0.address
		.servo_controllerv1_0_avalon_slave_0_write            (mm_interconnect_0_servo_controllerv1_0_avalon_slave_0_write),            //                                          .write
		.servo_controllerv1_0_avalon_slave_0_read             (mm_interconnect_0_servo_controllerv1_0_avalon_slave_0_read),             //                                          .read
		.servo_controllerv1_0_avalon_slave_0_readdata         (mm_interconnect_0_servo_controllerv1_0_avalon_slave_0_readdata),         //                                          .readdata
		.servo_controllerv1_0_avalon_slave_0_writedata        (mm_interconnect_0_servo_controllerv1_0_avalon_slave_0_writedata),        //                                          .writedata
		.sysid_qsys_control_slave_address                     (mm_interconnect_0_sysid_qsys_control_slave_address),                     //                  sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata                    (mm_interconnect_0_sysid_qsys_control_slave_readdata),                    //                                          .readdata
		.tc_instruct_mem_s2_address                           (mm_interconnect_0_tc_instruct_mem_s2_address),                           //                        tc_instruct_mem_s2.address
		.tc_instruct_mem_s2_write                             (mm_interconnect_0_tc_instruct_mem_s2_write),                             //                                          .write
		.tc_instruct_mem_s2_readdata                          (mm_interconnect_0_tc_instruct_mem_s2_readdata),                          //                                          .readdata
		.tc_instruct_mem_s2_writedata                         (mm_interconnect_0_tc_instruct_mem_s2_writedata),                         //                                          .writedata
		.tc_instruct_mem_s2_byteenable                        (mm_interconnect_0_tc_instruct_mem_s2_byteenable),                        //                                          .byteenable
		.tc_instruct_mem_s2_chipselect                        (mm_interconnect_0_tc_instruct_mem_s2_chipselect),                        //                                          .chipselect
		.tc_instruct_mem_s2_clken                             (mm_interconnect_0_tc_instruct_mem_s2_clken),                             //                                          .clken
		.timer_s1_address                                     (mm_interconnect_0_timer_s1_address),                                     //                                  timer_s1.address
		.timer_s1_write                                       (mm_interconnect_0_timer_s1_write),                                       //                                          .write
		.timer_s1_readdata                                    (mm_interconnect_0_timer_s1_readdata),                                    //                                          .readdata
		.timer_s1_writedata                                   (mm_interconnect_0_timer_s1_writedata),                                   //                                          .writedata
		.timer_s1_chipselect                                  (mm_interconnect_0_timer_s1_chipselect),                                  //                                          .chipselect
		.timestamp_s1_address                                 (mm_interconnect_0_timestamp_s1_address),                                 //                              timestamp_s1.address
		.timestamp_s1_write                                   (mm_interconnect_0_timestamp_s1_write),                                   //                                          .write
		.timestamp_s1_readdata                                (mm_interconnect_0_timestamp_s1_readdata),                                //                                          .readdata
		.timestamp_s1_writedata                               (mm_interconnect_0_timestamp_s1_writedata),                               //                                          .writedata
		.timestamp_s1_chipselect                              (mm_interconnect_0_timestamp_s1_chipselect),                              //                                          .chipselect
		.tmp101_s1_address                                    (mm_interconnect_0_tmp101_s1_address),                                    //                                 tmp101_s1.address
		.tmp101_s1_write                                      (mm_interconnect_0_tmp101_s1_write),                                      //                                          .write
		.tmp101_s1_read                                       (mm_interconnect_0_tmp101_s1_read),                                       //                                          .read
		.tmp101_s1_readdata                                   (mm_interconnect_0_tmp101_s1_readdata),                                   //                                          .readdata
		.tmp101_s1_writedata                                  (mm_interconnect_0_tmp101_s1_writedata),                                  //                                          .writedata
		.uart_rs485_s1_address                                (mm_interconnect_0_uart_rs485_s1_address),                                //                             uart_rs485_s1.address
		.uart_rs485_s1_write                                  (mm_interconnect_0_uart_rs485_s1_write),                                  //                                          .write
		.uart_rs485_s1_read                                   (mm_interconnect_0_uart_rs485_s1_read),                                   //                                          .read
		.uart_rs485_s1_readdata                               (mm_interconnect_0_uart_rs485_s1_readdata),                               //                                          .readdata
		.uart_rs485_s1_writedata                              (mm_interconnect_0_uart_rs485_s1_writedata)                               //                                          .writedata
	);

	DE0_CV_QSYS_mm_interconnect_1 mm_interconnect_1 (
		.pll_outclk0_clk                                          (pll_outclk0_clk),                                          //                                     pll_outclk0.clk
		.nios2_qsys_reset_reset_bridge_in_reset_reset             (rst_controller_001_reset_out_reset),                       //          nios2_qsys_reset_reset_bridge_in_reset.reset
		.nios2_qsys_tightly_coupled_instruction_master_0_address  (nios2_qsys_tightly_coupled_instruction_master_0_address),  // nios2_qsys_tightly_coupled_instruction_master_0.address
		.nios2_qsys_tightly_coupled_instruction_master_0_read     (nios2_qsys_tightly_coupled_instruction_master_0_read),     //                                                .read
		.nios2_qsys_tightly_coupled_instruction_master_0_readdata (nios2_qsys_tightly_coupled_instruction_master_0_readdata), //                                                .readdata
		.nios2_qsys_tightly_coupled_instruction_master_0_clken    (nios2_qsys_tightly_coupled_instruction_master_0_clken),    //                                                .clken
		.tc_instruct_mem_s1_address                               (mm_interconnect_1_tc_instruct_mem_s1_address),             //                              tc_instruct_mem_s1.address
		.tc_instruct_mem_s1_write                                 (mm_interconnect_1_tc_instruct_mem_s1_write),               //                                                .write
		.tc_instruct_mem_s1_readdata                              (mm_interconnect_1_tc_instruct_mem_s1_readdata),            //                                                .readdata
		.tc_instruct_mem_s1_writedata                             (mm_interconnect_1_tc_instruct_mem_s1_writedata),           //                                                .writedata
		.tc_instruct_mem_s1_byteenable                            (mm_interconnect_1_tc_instruct_mem_s1_byteenable),          //                                                .byteenable
		.tc_instruct_mem_s1_chipselect                            (mm_interconnect_1_tc_instruct_mem_s1_chipselect),          //                                                .chipselect
		.tc_instruct_mem_s1_clken                                 (mm_interconnect_1_tc_instruct_mem_s1_clken)                //                                                .clken
	);

	DE0_CV_QSYS_mm_interconnect_2 mm_interconnect_2 (
		.pll_outclk0_clk                                          (pll_outclk0_clk),                                          //                                     pll_outclk0.clk
		.boot_rom_reset1_reset_bridge_in_reset_reset              (rst_controller_reset_out_reset),                           //           boot_rom_reset1_reset_bridge_in_reset.reset
		.nios2_qsys_reset_reset_bridge_in_reset_reset             (rst_controller_001_reset_out_reset),                       //          nios2_qsys_reset_reset_bridge_in_reset.reset
		.nios2_qsys_tightly_coupled_instruction_master_1_address  (nios2_qsys_tightly_coupled_instruction_master_1_address),  // nios2_qsys_tightly_coupled_instruction_master_1.address
		.nios2_qsys_tightly_coupled_instruction_master_1_read     (nios2_qsys_tightly_coupled_instruction_master_1_read),     //                                                .read
		.nios2_qsys_tightly_coupled_instruction_master_1_readdata (nios2_qsys_tightly_coupled_instruction_master_1_readdata), //                                                .readdata
		.nios2_qsys_tightly_coupled_instruction_master_1_clken    (nios2_qsys_tightly_coupled_instruction_master_1_clken),    //                                                .clken
		.boot_rom_s1_address                                      (mm_interconnect_2_boot_rom_s1_address),                    //                                     boot_rom_s1.address
		.boot_rom_s1_write                                        (mm_interconnect_2_boot_rom_s1_write),                      //                                                .write
		.boot_rom_s1_readdata                                     (mm_interconnect_2_boot_rom_s1_readdata),                   //                                                .readdata
		.boot_rom_s1_writedata                                    (mm_interconnect_2_boot_rom_s1_writedata),                  //                                                .writedata
		.boot_rom_s1_byteenable                                   (mm_interconnect_2_boot_rom_s1_byteenable),                 //                                                .byteenable
		.boot_rom_s1_chipselect                                   (mm_interconnect_2_boot_rom_s1_chipselect),                 //                                                .chipselect
		.boot_rom_s1_clken                                        (mm_interconnect_2_boot_rom_s1_clken)                       //                                                .clken
	);

	DE0_CV_QSYS_irq_mapper irq_mapper (
		.clk           (pll_outclk0_clk),                    //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),           // receiver5.irq
		.sender_irq    (nios2_qsys_irq_irq)                  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (pll_outclk0_clk),                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_qsys_debug_reset_request_reset),   // reset_in1.reset
		.clk            (pll_outclk0_clk),                        //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
