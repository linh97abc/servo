module detect_hall_pos
(
    clk,
    reset_n,
    hall, // a, b, c
    position
)

input clk;
input reset_n;
input [2:0] hall;

output reg [31:0] position;

reg [2:0] hall_old;

wire [31:0] pos_next;
wire [31:0] pos_prev;

assign pos_next = position + 1'b1;
assign pos_prev = position - 1'b1;

always @(posedge clk) begin
    if (~reset_n) begin
        position <= 0;
        hall_old <= 0;
    end else begin
        hall_old <= hall;
        case ({hall, hall_old})
            {3'b001, 3'b101}: position <= pos_next;
            {3'b001, 3'b011}: position <= pos_prev;

            {3'b011, 3'b001}: position <= pos_next;
            {3'b011, 3'b010}: position <= pos_prev;

            {3'b010, 3'b011}: position <= pos_next;
            {3'b010, 3'b110}: position <= pos_prev;

            {3'b110, 3'b010}: position <= pos_next;
            {3'b110, 3'b100}: position <= pos_prev;

            {3'b100, 3'b110}: position <= pos_next;
            {3'b100, 3'b101}: position <= pos_prev;

            {3'b101, 3'b100}: position <= pos_next;
            {3'b101, 3'b001}: position <= pos_prev;

            default: position <= position;
        endcase
    end
end

endmodule